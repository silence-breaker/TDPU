`timescale 1ns / 1ps
package package_def;
  typedef enum logic [1:0] {
    W_ZERO = 2'b01,
    W_POS  = 2'b10,
    W_NEG  = 2'b00
  } weight_t;
endpackage
